
module addr_sel(Spc,Ssp);
input Spc,Ssp;


endmodule
