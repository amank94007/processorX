
module stack_ptr();


endmodule
