module alu_tb();
parameter ADD=1;
	parameter ADI=2;
	parameter ACA=3;
	parameter ACI=4;
	parameter SUB=5;
	parameter SCI=6;
	parameter SBI=7;
	parameter SCA=7;
	parameter XNR=9;
	parameter XNI=10;
	parameter XOR=11;
	parameter XRI=12;
	parameter AND=13;
	parameter ANI=14;
	parameter ORA=15;
	parameter ORI=16;
	parameter NOT=17;
	parameter NEG=18;
	parameter SRL=19;
	parameter SLL=20;
	parameter ASR=21;
	parameter ASL=22;
	parameter SRC=23;
	parameter SLC=24;
	parameter ROR=25;
	parameter ROL=26;
	parameter RRC=27;
	parameter RLC=28;
	parameter CLR=29;
	parameter INC=30;
	parameter DEC=31;
	parameter POP=32;
	parameter PSH=33;
	parameter MVS=34;
	parameter STS=35;
	parameter CCP=36;
	parameter JCP=37;
	parameter CCD=38;
	parameter JCD=39;
	parameter RTC=40;
	parameter JCA=41;
	parameter MVP=42;
	parameter RTU=43;
	parameter CUA=44;
	parameter STA=45;
	parameter CLA=46;
	parameter MVR=47;
	parameter JUA=48;
	parameter CUP=49;
	parameter JUP=50;
	parameter CUD=51;
	parameter JUD=52;
	parameter NOP=53;
wire [31:0]result;
wire [4:0]flags;
reg cin,fl,clkout;
reg [31:0]A,B,val;
reg [7:0]opcode;
alu a1(.result(result),.flags(flags),.A(A),.B(B),.opcode(opcode),.clkout(clkout),.cin(cin),.val(val),.fl(fl));
initial
clkout=0;
always
#5 clkout=~clkout;
initial
cin=0;fl=0;
#5  opcode=ADD;A=32'hABCD1234;B=32'hBCDABCAD;
#5	opcode=ADI;A=32'hABCD1235;
#5	opcode=ACA;A=32'hABCD1236;
#5	opcode=ACI;A=32'hABCD1237;
#5	opcode=SUB;A=32'hABCD1238;
#5	opcode=SCI;A=32'hABCD1239;
#5	opcode=SBI;A=32'hABCD123A;
#5	opcode=SCA;A=32'hABCD123B;
#5	opcode=XNR;A=32'hABCD123C;
#5	opcode=XNI;A=32'hABCD123D;
#5 opcode=XOR;A=32'hABCD123E;
#5 opcode=XRI;A=32'hABCD123F;
#5 opcode=AND;A=32'hABCD1240;
#5 opcode=ANI;A=32'hABCD1241;
#5 opcode=ORA;A=32'hABCD1234;
#5 opcode=ORI;A=32'hABCD1234;
#5 opcode=NOT;A=32'hABCD1234;
#5 opcode=NEG;A=32'hABCD1234;
#5 opcode=SRL;A=32'hABCD1234;
#5 opcode=SLL;A=32'hABCD1234;
#5 opcode=ASR;A=32'hABCD1234;
#5 opcode=ASL;A=32'hABCD1234;
#5 opcode=SRC;A=32'hABCD1234;
#5 opcode=SLC;A=32'hABCD1234;
#5 opcode=ROR;A=32'hABCD1234;
#5 opcode=ROL;A=32'hABCD1234;
#5 opcode=RRC;A=32'hABCD1234;
#5 opcode=RLC;A=32'hABCD1234;
#5 opcode=CLR;A=32'hABCD1234;
#5 opcode=INC;A=32'hABCD1234;
#5 opcode=DEC;A=32'hABCD1234;
#5 opcode=POP;A=32'hABCD1234;
#5 opcode=PSH;A=32'hABCD1234;
#5 opcode=MVS;A=32'hABCD1234;
#5 opcode=STS;A=32'hABCD1234;
#5 opcode=CCP;A=32'hABCD1234;
#5 opcode=JCP;A=32'hABCD1234;
#5 opcode=CCD;A=32'hABCD1234;
#5 opcode=JCD;A=32'hABCD1234;
#5 opcode=RTC;A=32'hABCD1234;
#5 opcode=JCA;A=32'hABCD1234;
#5 opcode=MVP;A=32'hABCD1234;
#5 opcode=RTU;A=32'hABCD1234;
#5 opcode=CUA;A=32'hABCD1234;
#5 opcode=STA;A=32'hABCD1234;
#5 opcode=CLA;A=32'hABCD1234;
#5 opcode=MVR;A=32'hABCD1234;
#5 opcode=JUA;A=32'hABCD1234;
#5 opcode=CUP;A=32'hABCD1234;
#5 opcode=JUP;A=32'hABCD1234;
#5 opcode=CUD;A=32'hABCD1234;
#5 opcode=JUD;A=32'hABCD1234;
#5 opcode=NOP;A=32'hABCD1234;